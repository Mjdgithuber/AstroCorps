<Level>
	<Size width="10" height="10"></Size>
	<Tile name="assets\blocks\tree.png" x="0" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="1" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="2" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="3" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="4" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="5" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="6" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="7" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="8" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="0"></Tile>
	<Tile name="assets\blocks\tree.png" x="0" y="1"></Tile>
	<Tile name="assets\blocks\z.png" x="1" y="1"></Tile>
	<Tile name="assets\blocks\grass.png" x="2" y="1"></Tile>
	<Tile name="assets\blocks\grass.png" x="3" y="1"></Tile>
	<Tile name="assets\blocks\grass.png" x="4" y="1"></Tile>
	<Tile name="assets\blocks\grass.png" x="5" y="1"></Tile>
	<Tile name="assets\blocks\grass.png" x="6" y="1"></Tile>
	<Tile name="assets\blocks\grass.png" x="7" y="1"></Tile>
	<Tile name="assets\blocks\grass.png" x="8" y="1"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="1"></Tile>
	<Tile name="assets\blocks\grass.png" x="0" y="2"></Tile>
	<Tile name="assets\blocks\grass.png" x="1" y="2"></Tile>
	<Tile name="assets\blocks\grass.png" x="2" y="2"></Tile>
	<Tile name="assets\blocks\grass.png" x="3" y="2"></Tile>
	<Tile name="assets\blocks\grass.png" x="4" y="2"></Tile>
	<Tile name="assets\blocks\grass.png" x="5" y="2"></Tile>
	<Tile name="assets\blocks\grass.png" x="6" y="2"></Tile>
	<Tile name="assets\blocks\grass.png" x="7" y="2"></Tile>
	<Tile name="assets\blocks\grass.png" x="8" y="2"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="2"></Tile>
	<Tile name="assets\blocks\tree.png" x="0" y="3"></Tile>
	<Tile name="assets\blocks\grass.png" x="1" y="3"></Tile>
	<Tile name="assets\blocks\grass.png" x="2" y="3"></Tile>
	<Tile name="assets\blocks\grass.png" x="3" y="3"></Tile>
	<Tile name="assets\blocks\z.png" x="4" y="3"></Tile>
	<Tile name="assets\blocks\grass.png" x="5" y="3"></Tile>
	<Tile name="assets\blocks\grass.png" x="6" y="3"></Tile>
	<Tile name="assets\blocks\grass.png" x="7" y="3"></Tile>
	<Tile name="assets\blocks\grass.png" x="8" y="3"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="3"></Tile>
	<Tile name="assets\blocks\tree.png" x="0" y="4"></Tile>
	<Tile name="assets\blocks\grass.png" x="1" y="4"></Tile>
	<Tile name="assets\blocks\grass.png" x="2" y="4"></Tile>
	<Tile name="assets\blocks\grass.png" x="3" y="4"></Tile>
	<Tile name="assets\blocks\grass.png" x="4" y="4"></Tile>
	<Tile name="assets\blocks\grass.png" x="5" y="4"></Tile>
	<Tile name="assets\blocks\grass.png" x="6" y="4"></Tile>
	<Tile name="assets\blocks\grass.png" x="7" y="4"></Tile>
	<Tile name="assets\blocks\grass.png" x="8" y="4"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="4"></Tile>
	<Tile name="assets\blocks\tree.png" x="0" y="5"></Tile>
	<Tile name="assets\blocks\grass.png" x="1" y="5"></Tile>
	<Tile name="assets\blocks\grass.png" x="2" y="5"></Tile>
	<Tile name="assets\blocks\grass.png" x="3" y="5"></Tile>
	<Tile name="assets\blocks\z.png" x="4" y="5"></Tile>
	<Tile name="assets\blocks\grass.png" x="5" y="5"></Tile>
	<Tile name="assets\blocks\grass.png" x="6" y="5"></Tile>
	<Tile name="assets\blocks\grass.png" x="7" y="5"></Tile>
	<Tile name="assets\blocks\grass.png" x="8" y="5"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="5"></Tile>
	<Tile name="assets\blocks\tree.png" x="0" y="6"></Tile>
	<Tile name="assets\blocks\grass.png" x="1" y="6"></Tile>
	<Tile name="assets\blocks\grass.png" x="2" y="6"></Tile>
	<Tile name="assets\blocks\grass.png" x="3" y="6"></Tile>
	<Tile name="assets\blocks\grass.png" x="4" y="6"></Tile>
	<Tile name="assets\blocks\grass.png" x="5" y="6"></Tile>
	<Tile name="assets\blocks\grass.png" x="6" y="6"></Tile>
	<Tile name="assets\blocks\grass.png" x="7" y="6"></Tile>
	<Tile name="assets\blocks\grass.png" x="8" y="6"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="6"></Tile>
	<Tile name="assets\blocks\tree.png" x="0" y="7"></Tile>
	<Tile name="assets\blocks\grass.png" x="1" y="7"></Tile>
	<Tile name="assets\blocks\grass.png" x="2" y="7"></Tile>
	<Tile name="assets\blocks\grass.png" x="3" y="7"></Tile>
	<Tile name="assets\blocks\grass.png" x="4" y="7"></Tile>
	<Tile name="assets\blocks\grass.png" x="5" y="7"></Tile>
	<Tile name="assets\blocks\grass.png" x="6" y="7"></Tile>
	<Tile name="assets\blocks\grass.png" x="7" y="7"></Tile>
	<Tile name="assets\blocks\grass.png" x="8" y="7"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="7"></Tile>
	<Tile name="assets\blocks\tree.png" x="0" y="8"></Tile>
	<Tile name="assets\blocks\grass.png" x="1" y="8"></Tile>
	<Tile name="assets\blocks\grass.png" x="2" y="8"></Tile>
	<Tile name="assets\blocks\grass.png" x="3" y="8"></Tile>
	<Tile name="assets\blocks\grass.png" x="4" y="8"></Tile>
	<Tile name="assets\blocks\grass.png" x="5" y="8"></Tile>
	<Tile name="assets\blocks\grass.png" x="6" y="8"></Tile>
	<Tile name="assets\blocks\grass.png" x="7" y="8"></Tile>
	<Tile name="assets\blocks\grass.png" x="8" y="8"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="8"></Tile>
	<Tile name="assets\blocks\tree.png" x="0" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="1" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="2" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="3" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="4" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="5" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="6" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="7" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="8" y="9"></Tile>
	<Tile name="assets\blocks\tree.png" x="9" y="9"></Tile>
</Level>
